module eightbit_alu(
	input[7:0] a, 
	input[7:0] b, 
	input[2:0] sel, 
	output reg[7:0] f,
	output reg ovf, 
	output reg take_branch);
	
	reg[8:0] a9, b9, f9;
	
	always @(a, b, sel)
	begin
		ovf = 0;
		take_branch = 0;
		case(sel)
			3'd0: 
			begin 
				a9 = a;
				b9 = b;
				f9 = a9 + b9;
				f = f9[7:0];
				ovf = f9[8];
			end
			3'd1:
				f = ~b;
			3'd2:
				f = a & b;
			3'd3:
				f = a | b;
			3'd4:
			begin 
				f[0] <= a[1];
				f[1] <= a[2];
				f[2] <= a[3];
				f[3] <= a[4];
				f[4] <= a[5];
				f[5] <= a[6];
				f[6] <= a[7];
				f[7] <= a[7];
			end
			3'd5:
			begin 
				f[0] <= 1'b0;
				f[1] <= a[0];
				f[2] <= a[1];
				f[3] <= a[2];
				f[4] <= a[3];
				f[5] <= a[4];
				f[6] <= a[5];
				f[7] <= a[6];
			end
			3'd6:
				take_branch = (a == b);
			3'd7:
				take_branch = (a != b);
		endcase
	end
endmodule

module Test;

	reg[7:0] a, b;
	reg[2:0] sel;
	wire[7:0] f;
	wire ovf, take_branch;

	eightbit_alu circuit(a, b, sel, f, ovf, take_branch);

	initial begin
		$monitor("%d a=%b b=%b sel=%d, f=%b overflow=%b branch=%b", 
			$time,
			a, b, sel, f, ovf, take_branch);

		#10 a = 0; b = 0; sel = 0;
		#10 a = 8'b00000000; b = 8'b11111111; sel = 0;
		#10 a = 8'b11111111; b = 8'b11111111; sel = 0;
		#10 a = 8'b10000000; b = 8'b10000000; sel = 0;
		#10 a = 8'b01000000; b = 8'b01000000; sel = 0;
		#10 a = 8'b00100000; b = 8'b00100000; sel = 0;
		#10 a = 8'b00010000; b = 8'b00010000; sel = 0;
		#10 a = 8'b00001000; b = 8'b00001000; sel = 0;
		#10 a = 8'b00000100; b = 8'b00000100; sel = 0;
		#10 a = 8'b00000010; b = 8'b00000010; sel = 0;
		#10 a = 8'b00000001; b = 8'b00000001; sel = 0;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 1;
		#10 a = 8'b00000000; b = 8'b11111111; sel = 1;
		#10 a = 8'b00000000; b = 8'b10101010; sel = 1;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 2;
		#10 a = 8'b11111111; b = 8'b00000000; sel = 2;
		#10 a = 8'b11111111; b = 8'b11111111; sel = 2;
		#10 a = 8'b10101010; b = 8'b10101010; sel = 2;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 3;
		#10 a = 8'b11111111; b = 8'b11111111; sel = 3;
		#10 a = 8'b11111111; b = 8'b00000000; sel = 3;
		#10 a = 8'b10101010; b = 8'b10101010; sel = 3;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 4;
		#10 a = 8'b00000001; b = 8'b00000000; sel = 4;
		#10 a = 8'b00000010; b = 8'b00000000; sel = 4;
		#10 a = 8'b00000100; b = 8'b00000000; sel = 4;
		#10 a = 8'b00001000; b = 8'b00000000; sel = 4;
		#10 a = 8'b00010000; b = 8'b00000000; sel = 4;
		#10 a = 8'b00100000; b = 8'b00000000; sel = 4;
		#10 a = 8'b01000000; b = 8'b00000000; sel = 4;
		#10 a = 8'b10000000; b = 8'b00000000; sel = 4;
		#10 a = 8'b11111111; b = 8'b00000000; sel = 4;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 5;
		#10 a = 8'b00000001; b = 8'b00000000; sel = 5;
		#10 a = 8'b00000010; b = 8'b00000000; sel = 5;
		#10 a = 8'b00000100; b = 8'b00000000; sel = 5;
		#10 a = 8'b00001000; b = 8'b00000000; sel = 5;
		#10 a = 8'b00010000; b = 8'b00000000; sel = 5;
		#10 a = 8'b00100000; b = 8'b00000000; sel = 5;
		#10 a = 8'b01000000; b = 8'b00000000; sel = 5;
		#10 a = 8'b10000000; b = 8'b00000000; sel = 5;
		#10 a = 8'b11111111; b = 8'b00000000; sel = 5;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 6;
		#10 a = 8'b11111111; b = 8'b11111111; sel = 6;
		#10 a = 8'b11111111; b = 8'b00000000; sel = 6;
		
		#10 a = 8'b00000000; b = 8'b00000000; sel = 7;
		#10 a = 8'b11111111; b = 8'b11111111; sel = 7;
		#10 a = 8'b11111111; b = 8'b00000000; sel = 7;
		
		#10 $finish; 

	end
endmodule
